module  bilinear_interpolation_rgb(


);





endmodule
