
// Efinity Top-level template
// Version: 2023.2.307.5.10
// Date: 2024-11-08 18:03

// Copyright (C) 2013 - 2023 Efinix Inc. All rights reserved.

// This file may be used as a starting point for Efinity synthesis top-level target.
// The port list here matches what is expected by Efinity constraint files generated
// by the Efinity Interface Designer.

// To use this:
//     #1)  Save this file with a different name to a different directory, where source files are kept.
//              Example: you may wish to save as C:\Users\Administrator\Desktop\wujisuofang\Ti60F225_ADV7611_HDMI_480P\Ti60_ADV7611_HDMI_640x480_EDID\Ti60_Demo.v
//     #2)  Add the newly saved file into Efinity project as design file
//     #3)  Edit the top level entity in Efinity project to:  Ti60_Demo
//     #4)  Insert design content.


module Ti60_Demo
(
  input clk_24m,
  input clk_25m,
  input cmos_ctl1,
  input [7:0] cmos_data,
  input cmos_href,
  input cmos_sdat_IN,
  input cmos_vsync,
  input sys_pll_lock,
  input ddr_pll_lock,
  input dsi_pll_lock,
  input lvds_pll_lock,
  input dsi_serclk_i,
  input dsi_txcclk_i,
  input dsi_refclk_i,
  input tdqss_clk,
  input tac_clk,
  input dsi_byteclk_i,
  input clk_pixel,
  input clk_sys,
  input clk_pixel_10x,
  input twd_clk,
  input csi_rxc_i,
  input clk_lvds_1x,
  input clk_27m,
  input core_clk,
  input clk_lvds_7x,
  input cmos_pclk,
  input clk_54m,
  input csi_ctl0_i,
  input csi_ctl1_i,
  input csi_scl_i,
  input csi_sda_i,
  input [15:0] i_dq_hi,
  input [15:0] i_dq_lo,
  input [1:0] i_dqs_hi,
  input [1:0] i_dqs_lo,
  input [1:0] i_dqs_n_hi,
  input [1:0] i_dqs_n_lo,
  input [23:0] hdmi_data_i,
  input hdmi_de_i,
  input hdmi_hs_i,
  input hdmi_pclk_i,
  input hdmi_sda_io_IN,
  input hdmi_vs_i,
  input uart_rx_i,
  input csi_rxc_lp_n_i,
  input csi_rxc_lp_p_i,
  input [7:0] csi_rxd0_hs_i,
  input csi_rxd0_lp_n_i,
  input csi_rxd0_lp_p_i,
  input [7:0] csi_rxd1_hs_i,
  input csi_rxd1_lp_n_i,
  input csi_rxd1_lp_p_i,
  input [7:0] csi_rxd2_hs_i,
  input csi_rxd2_lp_n_i,
  input csi_rxd2_lp_p_i,
  input [7:0] csi_rxd3_hs_i,
  input csi_rxd3_lp_n_i,
  input csi_rxd3_lp_p_i,
  input dsi_txd0_lp_n_i,
  input dsi_txd0_lp_p_i,
  input dsi_txd1_lp_n_i,
  input dsi_txd1_lp_p_i,
  input dsi_txd2_lp_n_i,
  input dsi_txd2_lp_p_i,
  input dsi_txd3_lp_n_i,
  input dsi_txd3_lp_p_i,
  output cmos_ctl2,
  output cmos_sclk,
  output cmos_sdat_OUT,
  output cmos_sdat_OE,
  output [5:0] led_o,
  output sys_pll_rstn_o,
  output ddr_pll_rstn_o,
  output [2:0] shift,
  output shift_ena,
  output [4:0] shift_sel,
  output dsi_pll_rstn_o,
  output lvds_pll_rstn_o,
  output hdmi_txc_oe,
  output [9:0] hdmi_txc_o,
  output hdmi_txc_rst_o,
  output hdmi_txd0_oe,
  output [9:0] hdmi_txd0_o,
  output hdmi_txd0_rst_o,
  output hdmi_txd1_oe,
  output [9:0] hdmi_txd1_o,
  output hdmi_txd1_rst_o,
  output hdmi_txd2_oe,
  output [9:0] hdmi_txd2_o,
  output hdmi_txd2_rst_o,
  output lvds_txc_oe,
  output [6:0] lvds_txc_o,
  output lvds_txc_rst_o,
  output lvds_txd0_oe,
  output [6:0] lvds_txd0_o,
  output lvds_txd0_rst_o,
  output lvds_txd1_oe,
  output [6:0] lvds_txd1_o,
  output lvds_txd1_rst_o,
  output lvds_txd2_oe,
  output [6:0] lvds_txd2_o,
  output lvds_txd2_rst_o,
  output lvds_txd3_oe,
  output [6:0] lvds_txd3_o,
  output lvds_txd3_rst_o,
  output [15:0] addr,
  output adv7611_rstn,
  output [2:0] ba,
  output cas,
  output cke,
  output clk_n_hi,
  output clk_n_lo,
  output clk_p_hi,
  output clk_p_lo,
  output cmos_ctl3,
  output cs,
  output csi_ctl0_o,
  output csi_ctl0_oe,
  output csi_ctl1_o,
  output csi_ctl1_oe,
  output csi_scl_o,
  output csi_scl_oe,
  output csi_sda_o,
  output csi_sda_oe,
  output [1:0] o_dm_hi,
  output [1:0] o_dm_lo,
  output [15:0] o_dq_hi,
  output [15:0] o_dq_lo,
  output [15:0] o_dq_oe,
  output [1:0] o_dqs_hi,
  output [1:0] o_dqs_lo,
  output [1:0] o_dqs_oe,
  output [1:0] o_dqs_n_hi,
  output [1:0] o_dqs_n_lo,
  output [1:0] o_dqs_n_oe,
  output dsi_pwm_o,
  output dsi_resetn_o,
  output hdmi_scl_io,
  output hdmi_sda_io_OUT,
  output hdmi_sda_io_OE,
  output odt,
  output ras,
  output reset,
  output spi_sck_o,
  output spi_ssn_o,
  output uart_tx_o,
  output we,
  output csi_rxc_hs_en_o,
  output csi_rxc_hs_term_en_o,
  output csi_rxd0_hs_en_o,
  output csi_rxd0_hs_term_en_o,
  output csi_rxd0_rst_o,
  output csi_rxd1_hs_en_o,
  output csi_rxd1_hs_term_en_o,
  output csi_rxd1_rst_o,
  output csi_rxd2_hs_en_o,
  output csi_rxd2_hs_term_en_o,
  output csi_rxd2_rst_o,
  output csi_rxd3_hs_en_o,
  output csi_rxd3_hs_term_en_o,
  output csi_rxd3_rst_o,
  output dsi_txc_hs_oe,
  output [7:0] dsi_txc_hs_o,
  output dsi_txc_lp_n_oe,
  output dsi_txc_lp_n_o,
  output dsi_txc_lp_p_oe,
  output dsi_txc_lp_p_o,
  output dsi_txc_rst_o,
  output dsi_txd0_hs_oe,
  output [7:0] dsi_txd0_hs_o,
  output dsi_txd0_lp_n_oe,
  output dsi_txd0_lp_n_o,
  output dsi_txd0_lp_p_oe,
  output dsi_txd0_lp_p_o,
  output dsi_txd0_rst_o,
  output dsi_txd1_hs_oe,
  output [7:0] dsi_txd1_hs_o,
  output dsi_txd1_lp_n_oe,
  output dsi_txd1_lp_n_o,
  output dsi_txd1_lp_p_oe,
  output dsi_txd1_lp_p_o,
  output dsi_txd1_rst_o,
  output dsi_txd2_hs_oe,
  output [7:0] dsi_txd2_hs_o,
  output dsi_txd2_lp_n_oe,
  output dsi_txd2_lp_n_o,
  output dsi_txd2_lp_p_oe,
  output dsi_txd2_lp_p_o,
  output dsi_txd2_rst_o,
  output dsi_txd3_hs_oe,
  output [7:0] dsi_txd3_hs_o,
  output dsi_txd3_lp_n_oe,
  output dsi_txd3_lp_n_o,
  output dsi_txd3_lp_p_oe,
  output dsi_txd3_lp_p_o,
  output dsi_txd3_rst_o
);


endmodule

